module tb ();
    
    initial begin
        $dumpfile("wave.vcd");
        $dumpvars;
    end

endmodule
